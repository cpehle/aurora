module descrambler(/*AUTOARG*/
   // Outputs
   descrambler_out,
   // Inputs
   clk, descrambler_in
   );
   input clk;
   input [63:0] descrambler_in;
   output [63:0] descrambler_out;


endmodule
