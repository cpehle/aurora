module aurora_descrambler(/*AUTOARG*/
   // Outputs
   aurora_descrambler_out,
   // Inputs
   aurora_descrambler_in
   );
   input [0:63] aurora_descrambler_in;
   output [0:63] aurora_descrambler_out;


endmodule
