module aurora_encoder();

endmodule
