module aurora_gearbox(/*AUTOARG*/);

endmodule
